--------------------------------------------------------------------------------
-- Entity:      Periferico_Copy
-- File:        Periferico_Copy.vhd
-- Description: DMA Controller for memory block transfer operations.
--              Handles bus arbitration (suspend) and data copy (memcpy).
-- Revision:    2.0 (Engineering Release)
-- Standard:    VHDL-93
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Periferico_Copy is
    Port ( 
        clock       : in  STD_LOGIC;
        reset       : in  STD_LOGIC;
        
        -- Bus Arbitration Interface
        suspend     : out STD_LOGIC; -- Request CPU Halt
        suspend_ack : in  STD_LOGIC; -- CPU Halted Acknowledge
        
        -- Master Memory Interface (Write-Only to System RAM)
        mem_address : out STD_LOGIC_VECTOR (31 downto 0);
        mem_data_out: out STD_LOGIC_VECTOR (31 downto 0);
        mem_we      : out STD_LOGIC; -- Write Enable (Active High)
        mem_ce      : out STD_LOGIC; -- Chip Enable
        mem_bw      : out STD_LOGIC; -- Byte Enable (1=Byte, 0=Word)
        
        -- Status Flag
        led_done    : out STD_LOGIC
    );
end Periferico_Copy;

architecture RTL of Periferico_Copy is

    -- FSM State Definitions
    type fsm_state_t is (
        ST_IDLE,        -- System Initialization
        ST_REQ_BUS,     -- Bus Request / Arbitration
        ST_FETCH_LAT,   -- Read Latency Wait State
        ST_TRANSFER,    -- Data Transfer Execution
        ST_PTR_INC,     -- Pointer Arithmetic
        ST_HALT         -- Operation Complete / Lock
    );
    
    signal current_state : fsm_state_t := ST_IDLE;

    -- Memory Pointers (Source and Destination)
    -- Base Source Address: 0x10012000 (Local ROM)
    signal ptr_read  : std_logic_vector(31 downto 0) := x"10012000";
    -- Base Dest Address:   0x10010020 (System RAM)
    signal ptr_write : std_logic_vector(31 downto 0) := x"10010020";
    
    -- Datapath Signals
    signal rom_clk_inv   : std_logic;
    signal rom_word_out  : std_logic_vector(31 downto 0);
    signal target_byte   : std_logic_vector(7 downto 0);

begin

    -- Clock Phase Inversion for Synchronous RAM
    rom_clk_inv <= not clock;

    -- =========================================================================
    -- LOCAL STORAGE INSTANTIATION (SOURCE DATA)
    -- =========================================================================
    -- NOTE: 'we' is hardwired to '1' to enforce READ-ONLY mode in the BRAM model
    -- generated by 'le_mars'. (Active Low Write Logic)
    SOURCE_MEMORY: entity work.data_mem_mod1 
    port map (
        clock       => rom_clk_inv, 
        ce          => '1',            
        we          => '1',            -- 1 = Read Mode / 0 = Write Mode
        bw          => '0',
        
        -- Address Decoding
        address     => ptr_read(12 downto 2),
        byte_choice => ptr_read(1 downto 0),
        
        data_in     => (others => '0'),
        data_out    => rom_word_out
    );

    -- =========================================================================
    -- BYTE STEERING LOGIC (Endianness Adjustment)
    -- =========================================================================
    -- Extracts the relevant byte from the 32-bit word based on address LSBs
    target_byte <= rom_word_out(7 downto 0)   when ptr_read(1 downto 0) = "00" else
                   rom_word_out(15 downto 8)  when ptr_read(1 downto 0) = "01" else
                   rom_word_out(23 downto 16) when ptr_read(1 downto 0) = "10" else
                   rom_word_out(31 downto 24);

    -- =========================================================================
    -- CONTROL FINITE STATE MACHINE (FSM)
    -- =========================================================================
    process(clock, reset)
    begin
        if reset = '1' then
            current_state <= ST_IDLE;
            -- Control Signals Reset
            suspend   <= '0';
            mem_we    <= '0'; mem_ce <= '0'; mem_bw <= '0';
            led_done  <= '0';
            -- Pointers Reset
            ptr_read  <= x"10012000";
            ptr_write <= x"10010020";
            
        elsif rising_edge(clock) then
            case current_state is
                
                -- State: System Idle / Reset Release
                when ST_IDLE =>
                    suspend <= '1'; -- Assert Bus Request
                    if suspend_ack = '1' then
                        current_state <= ST_FETCH_LAT;
                    else
                        current_state <= ST_IDLE;
                    end if;

                -- State: Memory Read Latency
                when ST_FETCH_LAT =>
                    -- Wait 1 cycle for BRAM output stabilization
                    mem_we <= '0';
                    mem_ce <= '0';
                    current_state <= ST_TRANSFER;

                -- State: Data Write to System RAM
                when ST_TRANSFER =>
                    mem_address <= ptr_write;
                    
                    -- Byte Replication for 32-bit Bus Alignment
                    mem_data_out <= target_byte & target_byte & target_byte & target_byte;
                    
                    mem_ce <= '1'; 
                    mem_we <= '1'; 
                    mem_bw <= '1'; -- Byte-Write Mode

                    -- Null Terminator Check (End of String)
                    if target_byte = x"00" then
                        current_state <= ST_HALT;
                    else
                        current_state <= ST_PTR_INC;
                    end if;

                -- State: Address Pointer Increment
                when ST_PTR_INC =>
                    mem_we <= '0';
                    mem_ce <= '0';
                    ptr_read  <= ptr_read + 1;
                    ptr_write <= ptr_write + 1;
                    current_state <= ST_FETCH_LAT;

                -- State: Operation Completed
                when ST_HALT =>
                    mem_we    <= '0';
                    mem_ce    <= '0';
                    suspend   <= '0';  -- Release Bus Control
                    led_done  <= '1';  -- Signal Completion
                    current_state <= ST_HALT; -- Lock State
                    
                when others =>
                    current_state <= ST_IDLE;
            end case;
        end if;
    end process;

end RTL;