--
--  Automatically Generated--  Authors: Fernando Moraes & Ney Calazans
--  Generation date: Tue Dec 09 14:06:44 2025
--

--------------------------------------------------------
--  Instruction Memory Module 1
--    512 32-bit words (2KBytes, 16Kbits, 1 BRAM)
--------------------------------------------------------
library IEEE;
use IEEE.Std_Logic_1164.all;
library UNISIM;
use UNISIM.vcomponents.all; 

entity program_memory is
    port( clock: in std_logic;
          address: in std_logic_vector(8 downto 0);
          instruction: out std_logic_vector(31 downto 0));
end program_memory;

architecture program_memory of program_memory is     
begin
           
   inst_mem : RAMB16_S36
   generic map (
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000008100000",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
            CLK     => clock,
            ADDR    => address,
            EN      => '1',
            WE      => '0',
            DI      => x"00000000",
            DIP     => x"0",
            DO      => instruction,
            SSR     => '0'
            );

end program_memory;

----------------------------------------------------------
--  Data Memory Module 0 - Four 2048 8-bit bytes blocks,
--      interleaved (8KBytes, 64Kbits, 4 BRAMs)
--  This module start address is 0x10010000
--  Possible data access methods for read/write operations:
--      * byte, at any address
--      * 32-bit words at addresses multiple of 4
--  When using more than one Memory Module beware:
--      1) Modules are independent of each other,
--          i.e. external decoding will define their
--          relative position in the memory map
--      2) Modules have 13-bit address lines in the
--          range 0x0000 - 0x1FFF. The most significant
--          11 bits are the signal named address. The 2
--          least significant bits are signal byte_choice.
--          In fact, the latter specify in which memory
--          block resides the byte in byte access. For
--          word access, byte_choice must be 00.
--
--  Interleaved memory Example: A memory with contents:
--  00 00 00 00
--  10 00 00 AA
--  20 00 BB 00
--  30 CC 00 00
--  
--  Will result in BRAM data memory first lines filled as:
--  
-- mem 3-  INIT_00 => X"...000000000000000000030201000",
-- mem 2-  INIT_00 => X"...0000000000000000000CC000000",
-- mem 1-  INIT_00 => X"...000000000000000000000BB0000",
-- mem 0-  INIT_00 => X"...00000000000000000000000AA00",
--
----------------------------------------------------------
library IEEE;
use IEEE.Std_Logic_1164.all;
library UNISIM;
use UNISIM.vcomponents.all; 

entity data_mem_mod0 is
    port( clock, ce, -- For now, ce is unused in module,
    	             -- The EN input of all blocks is '1'.
          we, bw: in std_logic;
          address: in std_logic_vector(10 downto 0);    -- 11 bits - 2048 addressable words
          byte_choice: in std_logic_vector(1 downto 0); -- 2 bits  - 1 of 4 addressable bytes
          data_in: in std_logic_vector(31 downto 0);
          data_out: out std_logic_vector(31 downto 0));
end data_mem_mod0;

architecture data_mem_mod0 of data_mem_mod0 is 
    signal we3, we2, we1, we0 : std_logic;
    signal d_in_mem3, d_in_mem2, d_in_mem1, d_in_mem0 : std_logic_vector(7 downto 0);
begin

    we3 <= '1' when (we='0' and ((bw='0') or (bw='1' and byte_choice="11"))) else '0';
    we2 <= '1' when (we='0' and ((bw='0') or (bw='1' and byte_choice="10"))) else '0';
    we1 <= '1' when (we='0' and ((bw='0') or (bw='1' and byte_choice="01"))) else '0';
    we0 <= '1' when (we='0' and ((bw='0') or (bw='1' and byte_choice="00"))) else '0';
    d_in_mem3 <= data_in(7 downto 0) when bw='1' else data_in(31 downto 24);
    d_in_mem2 <= data_in(7 downto 0) when bw='1' else data_in(23 downto 16);
    d_in_mem1 <= data_in(7 downto 0) when bw='1' else data_in(15 downto 8);
    d_in_mem0 <= data_in(7 downto 0);

   ----------------------------------------------------------------------------------
   -- bytes 31 a 24
   ----------------------------------------------------------------------------------
    block_3: RAMB16_S9
         generic map (
        INIT_00 => X"0000000000000000000000000000000000000000000000000074356374747565",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
         CLK     => clock,
         ADDR    => address,
         EN      => '1',
         WE      => we3,
         DI      => d_in_mem3,
         DIP     => "0",
         DO      => data_out(31 downto 24),
         SSR     => '0'
         );

   ----------------------------------------------------------------------------------
   -- bytes 23 a 16
   ----------------------------------------------------------------------------------
    block_2: RAMB16_S9
         generic map (
        INIT_00 => X"0000000000000000000000000000000000000000000000000078655363654a6d",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
         CLK     => clock,
         ADDR    => address,
         EN      => '1',
         WE      => we2,
         DI      => d_in_mem2,
         DIP     => "0",
         DO      => data_out(23 downto 16),
         SSR     => '0'
         );

   ----------------------------------------------------------------------------------
   -- bytes 15 a 8
   ----------------------------------------------------------------------------------
    block_1: RAMB16_S9
         generic map (
        INIT_00 => X"00000000000000000000000000000000000000000000000000746e2d4169266f",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
         CLK     => clock,
         ADDR    => address,
         EN      => '1',
         WE      => we1,
         DI      => d_in_mem1,
         DIP     => "0",
         DO      => data_out(15 downto 8),
         SSR     => '0'
         );

   ----------------------------------------------------------------------------------
   -- bytes 7 a 0
   ----------------------------------------------------------------------------------
    block_0: RAMB16_S9
         generic map (
        INIT_00 => X"000000000000000000000000000000000000000000000000002e65315f6c6f52",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
         CLK     => clock,
         ADDR    => address,
         EN      => '1',
         WE      => we0,
         DI      => d_in_mem0,
         DIP     => "0",
         DO      => data_out(7 downto 0),
         SSR     => '0'
         );

end data_mem_mod0;

----------------------------------------------------------
--  Data Memory Module 1 - Four 2048 8-bit bytes blocks,
--      interleaved (8KBytes, 64Kbits, 4 BRAMs)
--  This module start address is 0x10012000
--  Possible data access methods for read/write operations:
--      * byte, at any address
--      * 32-bit words at addresses multiple of 4
--  When using more than one Memory Module beware:
--      1) Modules are independent of each other,
--          i.e. external decoding will define their
--          relative position in the memory map
--      2) Modules have 13-bit address lines in the
--          range 0x0000 - 0x1FFF. The most significant
--          11 bits are the signal named address. The 2
--          least significant bits are signal byte_choice.
--          In fact, the latter specify in which memory
--          block resides the byte in byte access. For
--          word access, byte_choice must be 00.
--
--  Interleaved memory Example: A memory with contents:
--  00 00 00 00
--  10 00 00 AA
--  20 00 BB 00
--  30 CC 00 00
--  
--  Will result in BRAM data memory first lines filled as:
--  
-- mem 3-  INIT_00 => X"...000000000000000000030201000",
-- mem 2-  INIT_00 => X"...0000000000000000000CC000000",
-- mem 1-  INIT_00 => X"...000000000000000000000BB0000",
-- mem 0-  INIT_00 => X"...00000000000000000000000AA00",
--
----------------------------------------------------------
library IEEE;
use IEEE.Std_Logic_1164.all;
library UNISIM;
use UNISIM.vcomponents.all; 

entity data_mem_mod1 is
    port( clock, ce, -- For now, ce is unused in module,
    	             -- The EN input of all blocks is '1'.
          we, bw: in std_logic;
          address: in std_logic_vector(10 downto 0);    -- 11 bits - 2048 addressable words
          byte_choice: in std_logic_vector(1 downto 0); -- 2 bits  - 1 of 4 addressable bytes
          data_in: in std_logic_vector(31 downto 0);
          data_out: out std_logic_vector(31 downto 0));
end data_mem_mod1;

architecture data_mem_mod1 of data_mem_mod1 is 
    signal we3, we2, we1, we0 : std_logic;
    signal d_in_mem3, d_in_mem2, d_in_mem1, d_in_mem0 : std_logic_vector(7 downto 0);
begin

    we3 <= '1' when (we='0' and ((bw='0') or (bw='1' and byte_choice="11"))) else '0';
    we2 <= '1' when (we='0' and ((bw='0') or (bw='1' and byte_choice="10"))) else '0';
    we1 <= '1' when (we='0' and ((bw='0') or (bw='1' and byte_choice="01"))) else '0';
    we0 <= '1' when (we='0' and ((bw='0') or (bw='1' and byte_choice="00"))) else '0';
    d_in_mem3 <= data_in(7 downto 0) when bw='1' else data_in(31 downto 24);
    d_in_mem2 <= data_in(7 downto 0) when bw='1' else data_in(23 downto 16);
    d_in_mem1 <= data_in(7 downto 0) when bw='1' else data_in(15 downto 8);
    d_in_mem0 <= data_in(7 downto 0);

   ----------------------------------------------------------------------------------
   -- bytes 31 a 24
   ----------------------------------------------------------------------------------
    block_3: RAMB16_S9
         generic map (
        INIT_00 => X"6e6c65616e6f997220475254460d6e617468666f6569530a6553200a74756e65",
        INIT_01 => X"776f6f200a6c61736e6420574d5620430d726e0a65634865656169657920740a",
        INIT_02 => X"206f68656573746e20207777414953520d67746f20992c0a686e65642c619965",
        INIT_03 => X"6447736e656570746c6d76750a20616e6320657065762c746f2e6c68746f6462",
        INIT_04 => X"0d666c2020206f65754e4e45530a2e65792c4e4e45520a21746479742e4e616e",
        INIT_05 => X"616965732072436f65746165626e204e4e45520a2e6d207268696f687361666b",
        INIT_06 => X"746d6c676e746774616c7320202075206e0d22737679226c6b0d69656c74616c",
        INIT_07 => X"74646155657274616173616e6c676d6554500d2e6b207465642c6f4269722c6f",
        INIT_08 => X"49682c69736d6868656420646e696c756663207374202c0d797474206c6c206f",
        INIT_09 => X"74756472766e2068740a64746576496574206f57770d206e6f202e6f742c776c",
        INIT_0A => X"676d65726f2e6774206f69e26e7380656c6c20680a619964722069616e70770d",
        INIT_0B => X"6f746c6f20722c7420206f762c682c680d6320746161634d790a6e69206f6e6c",
        INIT_0C => X"776d7473666b6e692c722c0d6f6f77206d2020696863714170657474756e736e",
        INIT_0D => X"737961632020e2206c48732063202070616475720d6c4373206769792c204e2e",
        INIT_0E => X"6e742075736e74206d610d550a2e6574746472204e4f9945410a736120572020",
        INIT_0F => X"207461722065646520536c20736c75616f6e650a6963666175686320990d7573",
        INIT_10 => X"2074796945410a747420200a6972652020206f69e27273804e4f9945410a656d",
        INIT_11 => X"6f4f6e65686e746877689964740a6169536f4f520d61616f642075616f693f74",
        INIT_12 => X"656e2061686d200d672062206320206574652c4f520d736f6f494d560a3f6972",
        INIT_13 => X"7276797373730a616f684566736f636f79659461996f45206c6a69200d696f65",
        INIT_14 => X"656e752c0a6166632020616c496e6561650d6f736c7272e264726f4177207769",
        INIT_15 => X"2e69696c206165202080206f2c697461723f20746f7220640d616479a8656520",
        INIT_16 => X"68204376202061740a7365612e20692065630a657420627520697379730a410a",
        INIT_17 => X"20646869200d6b207268616f6579770d696c72747220206c5463636120777263",
        INIT_18 => X"0a6f75657420696865554c540d2020747272206d6b6f6f790d550a2e206f696f",
        INIT_19 => X"6569e2410a3f7365206f54500d746e68746520206e730a696e6d726969686969",
        INIT_1A => X"747320416e6c6774206b6d73620a6e202020637420686e6f54500d6f52617668",
        INIT_1B => X"6f6d2048777320206865686f6f6c202e6f65766c202075766554696f61616568",
        INIT_1C => X"726961682c7020742068686c2073496d66746f6b2e6920656554746561646820",
        INIT_1D => X"e22e75206e6c61756573200d420d746672656c7369736c6e2c6f65746f70616e",
        INIT_1E => X"6f757272726168200d202e6868733f206420682e75206c7320550a2e2064746c",
        INIT_1F => X"80796f616f656c750d7320676169206b6ce20a75796e6c73476972656e996f2e",
        INIT_20 => X"74683f646f997379797365750d202c6f45410a6d2069e26c20574c540d6d7420",
        INIT_21 => X"6f7220202072202c7365946d7380794d6d616f73750d686f496f68732061796b",
        INIT_22 => X"706e6154590a7468207263612e756f6b6ce22c686f746c6f746c6f7274710a67",
        INIT_23 => X"686f7220746261746c202e746765667274206d206c6d6b0d74206f6c6c68206f",
        INIT_24 => X"6f20682066204922688069206b204f0a7365226c20727420746e2c776e656f2c",
        INIT_25 => X"68747574206f6f6473612c7270696c7773200d68697374202069206868642069",
        INIT_26 => X"6e200a696e772074647261630a636f6420796f6f6f6d6c640a490a2e6b642074",
        INIT_27 => X"6f6e73206974650a4d0d7320736c79206d206d200a63207368e2727068642068",
        INIT_28 => X"2061616f70742c61612c740d4f0a657020206d68617320727041454a0d746570",
        INIT_29 => X"450a2e73e279202072677476746f7453454a0d61642074697420686e2072650d",
        INIT_2A => X"0d4c0d6475697320697973206d20542e2073650d6120667372726d6974652054",
        INIT_2B => X"222e67696d204764757473617220696d72694f520d6f767920747374696d6165",
        INIT_2C => X"72646f65206c0a6f7464206563682079610a520d6b206862696f454a0d65656b",
        INIT_2D => X"206e792067640d756566646573656d4872682072454e0d682020740a4d0d2e74",
        INIT_2E => X"6b6374616c0a6820686c6368686f6c496c696574796865757264750a75726465",
        INIT_2F => X"2e672c41494e0d7420e220736679746372203f752068496561450a2e6176654e",
        INIT_30 => X"0a6e65746e61706574204e45410a73752065202065202c0d4f0a736574696f65",
        INIT_31 => X"6e6f6e6c6765207961496c756b742c7457739920732072747562696669722068",
        INIT_32 => X"4a62412e72206ce22e6c78747979626173412e2073742c742043727372650a74",
        INIT_33 => X"62646669646e650d550a6174207920577320682043454a0d696f692075686e65",
        INIT_34 => X"e257454a0d68746779206949612c61454e0d6f6f6f69736f616599610d4c0d6f",
        INIT_35 => X"c36162202e6772652e6e68610a490a2e206b454e0d6e7464776865206c207420",
        INIT_36 => X"61207920206f546574206e6f52206e48226e65454e0d626977206f6b7376200d",
        INIT_37 => X"76667420696f0d616f7720206f75656c200a7479206d207265206f0a490a2e6e",
        INIT_38 => X"0a6e7665652068204c0d7320e2576973740a520d7965c36f206c7520546d2074",
        INIT_39 => X"680d6f726c72612020779965650a6f2c41530a2e6c2e6820616e0d68206e496f",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000002e65",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
         CLK     => clock,
         ADDR    => address,
         EN      => '1',
         WE      => we3,
         DI      => d_in_mem3,
         DIP     => "0",
         DO      => data_out(31 downto 24),
         SSR     => '0'
         );

   ----------------------------------------------------------------------------------
   -- bytes 23 a 16
   ----------------------------------------------------------------------------------
    block_2: RAMB16_S9
         generic map (
        INIT_00 => X"20656868615080654e4e45530a22696e697420636d76220d6e20740d654a616d",
        INIT_01 => X"7420206c0d206872616f6e20475244450a65650d70732068722068486165200d",
        INIT_02 => X"74637476726c7369656820414d5620490a6e206673806f0d7375686e7368806d",
        INIT_03 => X"6e2075696c74202020206f6f0d2c2061726663206d61752047657074206c7270",
        INIT_04 => X"2c206c6472646f726f414953520d79726f79414953490d6e6f6e6e6e6c200a6f",
        INIT_05 => X"207242792c650a6f72202068206e65414953490d726174677420666720202073",
        INIT_06 => X"206f740a61732020206f757364747072450a65616f65206161726c6720202069",
        INIT_07 => X"69656c0a6f69206868654c6574206f5745410a7373726f686e6f762074656f52",
        INIT_08 => X"20537961652074536320792020576c6f6f692c737379682e0a697561616c7363",
        INIT_09 => X"206f6e6f20726520610d20207361206d6e2c630a6f757220636d736361727399",
        INIT_0A => X"206f7761596520992c6774206f69e273707573630d658061696120746973206c",
        INIT_0B => X"7968204d2e69746f642172696c206c20226e7920206c6922610d61732c436574",
        INIT_0C => X"206f72202d6f75686869682068746f736f653b66746e200a756c20207461656b",
        INIT_0D => X"72206c6e77742067200a79676e727420206e6f6f2c75207564207361742c0a6c",
        INIT_0E => X"20992c6d2020992c206854500d737972206199794943804c430d6120650a6466",
        INIT_0F => X"6e20206179776e76650a6c74616b712063656d0d74756f696e746e73802e6d20",
        INIT_10 => X"6c2020574c430d72206e730d7365206e732e6d74206f69e24943804c430d6b20",
        INIT_11 => X"790a616863656f6320748061610d6d762074450a2e2065777261627773487420",
        INIT_12 => X"686f736873657421696e2073726568746f684f450a2e206e6e2047520d746e65",
        INIT_13 => X"746f772077200d656f7420207566696f744280658069206e65207273746e2068",
        INIT_14 => X"68696f640d746f6172687799206f7265682e68776565656f6165790a6f682070",
        INIT_15 => X"746e686c7965757772e24946747369656f776c206c6179692e68756dc36c6b2c",
        INIT_16 => X"74650a61657364610d742050792c70796d740d756e61206f2c6f6962690d420d",
        INIT_17 => X"642020726f2c20666f20207468626f3f6e6f75616f6472660a61692068206520",
        INIT_18 => X"0d666f756e6120746c0a410a3f756d736f653f73206e686854500d6e616e2068",
        INIT_19 => X"685420420d74696d675945410a682074696c727472200d70696f656820746176",
        INIT_1A => X"20202c0a6174207261696972200d6f6d742e206e2c74654345410a65206c2074",
        INIT_1B => X"6820650a6f696c66747774666e754968796e6f6c64737420620a6820726e5674",
        INIT_1C => X"70612053747375206877746c79690a696f6f6e6174746572720a6e6770202065",
        INIT_1D => X"497467736969207368747454590a73206f6362206d656c417372732020202065",
        INIT_1E => X"476f6f65656d746d2e6f6c732020796e6f2c576464656c2054500d6d656e6f6c",
        INIT_1F => X"e2206f2d6373696f2c65796e207461616c750d6f6d656c20206875202080596f",
        INIT_20 => X"2054646e7380496f6320726f2e6f6f474c430d61617420632c0a410a2120206c",
        INIT_21 => X"637065752e6179642057806969e27220207263756f2e776e2079742065686163",
        INIT_22 => X"2065504c540d72202c652068747179616c4965736668206d68204d6f65200d20",
        INIT_23 => X"73697473202072696c4967652072696920656568662061676572687569746566",
        INIT_24 => X"777974656f490a6420e26c67614f520d74200a6c7499746f726f747369734e6c",
        INIT_25 => X"63206f61686d546e206573672068627470793a7420206e652c727920546e7468",
        INIT_26 => X"69720d68696f6e6f20656d690d756f6e722072647969696f0d4c0d73206e6169",
        INIT_27 => X"68617073616f760d4f0a739972616c736c6f6c640d756f6420736720746e6520",
        INIT_28 => X"7368686469657473656e204f520d79206574207468702c67200a490a3f206d20",
        INIT_29 => X"4d0d6520736172746775206f6f646e0a490a2e70206e2061732c74613a70682e",
        INIT_2A => X"54550a657020202c686270796f730a727369482e74746699657020686f766e0a",
        INIT_2B => X"0a6e617320650a6520652070743f6c206653450a2e746165742020206c206868",
        INIT_2C => X"6572747674750d796972617620747220640d550a6f9974206b59490a22687320",
        INIT_2D => X"61616464206e2c6f686f61686968200a6f632c61530a3f747273610d4f0a726f",
        INIT_2E => X"6e202068610d2064202020742079650a61776b202074746165656e0d6f696e73",
        INIT_2F => X"6565790a4c450a6273657969694d6e63614f747061732064224d0d79206f7320",
        INIT_30 => X"0d6f62202070206d6e2c0a4c430d65207372652e666f794f520d656861207068",
        INIT_31 => X"20476574206e2c20680a6c6f6e206e2020208074492e612071206c206c746520",
        INIT_32 => X"20202274206f6c4965206169616d2072200a646f99656e20652065656f720d68",
        INIT_33 => X"696c6f656e6f68454e0d6d6e64207420722c74650a490a22787467654e746169",
        INIT_34 => X"740a490a2e63656e202c682068794d530a3f6420206f696e6868806854550a69",
        INIT_35 => X"696d206673207568652020200d4c0d747720530a3f616f6c207472736c742073",
        INIT_36 => X"6572206e79200a756e6161652065200a677272530a2e2064206574696961792c",
        INIT_37 => X"6f6f72736772216c746f642c6e2073726f0d616c796f67707679200d4c0d7965",
        INIT_38 => X"0d20656e6c657254550a697374206899610d550a6d20686c65206d740a207369",
        INIT_39 => X"542e6761616572652e61806c6d0d6e6e20520d7475227473634f2e7464612020",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000007420",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
         CLK     => clock,
         ADDR    => address,
         EN      => '1',
         WE      => we2,
         DI      => d_in_mem2,
         DIP     => "0",
         DO      => data_out(23 downto 16),
         SSR     => '0'
         );

   ----------------------------------------------------------------------------------
   -- bytes 15 a 8
   ----------------------------------------------------------------------------------
    block_1: RAMB16_S9
         generic map (
        INIT_00 => X"736820747020e268414953520d2e6b207772652067720a35652c630a6920206f",
        INIT_01 => X"20656e6c656c73656d6f654e4e454e530d68726161203f6374747320776b6f74",
        INIT_02 => X"72200a6f206f206f68747920475254460d696c2069e26f64612074616420e220",
        INIT_03 => X"696e5320207265742c736c6873642c70616f656120736f640a7420206b206175",
        INIT_04 => X"7264616e6f656c61594d5620490a642062414d5620480a6150616f416c640d74",
        INIT_05 => X"6b62206f79650d74656465207461574d5620480a65686120202c207564726461",
        INIT_06 => X"6e776e0d2065656c2c686f696e656165220d64206d682e207465206e65642c68",
        INIT_07 => X"7775700d746565207469206d6e2c630a4c430d7261650a7461696e2c754d6520",
        INIT_08 => X"2c0a74646b7420206e6f6e776c0a617920687365696d41750d776f2077696e20",
        INIT_09 => X"64636173616f76496879656e20682e6565656c0d6e6f616520416e2068612080",
        INIT_0A => X"2c6320200a6e73806520992c67542061206f61752c20e26c612065207269416c",
        INIT_0B => X"2067650a7367696f6e6d20676c616c412e616564737073206c2c697565206d6e",
        INIT_0C => X"73636f72646f20746173412e202072696f6865202065640d2062656e20207620",
        INIT_0D => X"757420696f99736e770d616e617573654961794674706e6f6f2c206e69790d6c",
        INIT_0E => X"738068207473806e2c5745410a7220692c4c80425320e2550a3f6d6e720d6e6c",
        INIT_0F => X"65642c65747461696d0d69692063207465506f2c6e4c207420206969e2682074",
        INIT_10 => X"6c756c20550a2e69736f692e2064736f696520992c6d540a5320e2550a2e7365",
        INIT_11 => X"200d6874692064697420e26c6822677261224d0d6f73797461202020200a6165",
        INIT_12 => X"747067202065497472726f656f68632064730a4d0d722c206b4e4e450a686b64",
        INIT_13 => X"20646f616f6f2e647472722c20207274750ae220e2686e697768204168206b63",
        INIT_14 => X"2068746e6473206c656320802c64756d5473736f666899206c64200d7274676f",
        INIT_15 => X"68207469746272616565200a68202077466f6c6520656d446420722073626173",
        INIT_16 => X"696d0d6c68652068226965226f72616d206520676f206468657668206854590a",
        INIT_17 => X"616d6574546e796f6e646b7374204e796d736f20636e65200d66746e74647672",
        INIT_18 => X"2c2020676f207320630d420d6f6f722066686e6e2c20205745410a6920206420",
        INIT_19 => X"209954590a69206f6e0a4c430d6773206e6f75616f6f65732063682074206c20",
        INIT_1A => X"796f640d6d6e796f206c6861652e6c69657a65656520740a4c430d6d6e6c7420",
        INIT_1B => X"206e720d74686c6f6c202020206f0a74207267656e757261200d2073626f2075",
        INIT_1C => X"2066770a63656f66632020696d200d68206e20546e61626f650d6561736d6f73",
        INIT_1D => X"0a732069617668207769494c540d6161666e6d676562690a6e66656674646573",
        INIT_1E => X"20792068742020416f476c2079496f616f740a656e62616545410a6972656e99",
        INIT_1F => X"752c686b2020775973756d6f7975206d996f2c73206d6164212064746ce20a74",
        INIT_20 => X"730a656920e22062756161596f677420550a2e6820992c6e790d420d6e65656c",
        INIT_21 => X"6e20726f73656d696c0ae2747420722e7974206d5974206b2e20616f63636d69",
        INIT_22 => X"65690a410a21617979652c576520206d990a6d20206765206765202069652e2c",
        INIT_23 => X"20736e69742c6477690a6e65746564656e6c727320734d6e6565636677696372",
        INIT_24 => X"6e6d696e72200d6e7374756e74450a2269650d6173806974656365206d200a6c",
        INIT_25 => X"7568726874730a6179726d6c67732020694d73206e65656865686c730a617374",
        INIT_26 => X"616f3b7420686f76796e20682c6d7461756777202072706f54550a7372652077",
        INIT_27 => X"20206974736e614f520d698065706f696174616e2c6f646e996d6c7420617673",
        INIT_28 => X"642077206c6c6e2064654f450a2e616e7373792074696d6c2c0d4c0d6f736c79",
        INIT_29 => X"4f0a6b9972726f6e206f2c6d6e20690d4c0d72736f726866657520727920546f",
        INIT_2A => X"454a0d67206e79657420696d72750d65656b226520636580792065776e6f650d",
        INIT_2B => X"0d69202065760d67796573732073206d200a4d0d6b206868616e657320652054",
        INIT_2C => X"6861206f654a2e20776f2061726f752c61454e0d6f80207320204c0d2e207365",
        INIT_2D => X"2020616f6141656874206c742074720d6c61794d520d726f6569684f520d656d",
        INIT_2E => X"696565206872666c796e74202c20740d68206c75742068646873202e75766169",
        INIT_2F => X"6e62610d4f420d65996f6d206c207561650a656120202069204f0a61736d722e",
        INIT_30 => X"2e67207465652c6565790d550a2e7279696f6872207341450a2e627420747354",
        INIT_31 => X"64206d6e746f756b740d6179614965793f6ee2690a7377746e686f6766207665",
        INIT_32 => X"746c0a737974990a7473772066202c722c0d6574806c656e6d2e6868746f2067",
        INIT_33 => X"546f2068617354530a3f65656e73612e7572696d0d4c0d2e652065732020206c",
        INIT_34 => X"610d4c0d6f755075656b742c74720a520d722074676720207420e257454a0d72",
        INIT_35 => X"7220654965654e546d736b6f54550a6f6f49520d65646e75742065776f616599",
        INIT_36 => X"7275666f6c650d676f20206d736d730d6e7522520d6467647962206c20724d64",
        INIT_37 => X"6c20697569506520206e6e6e6b6e20616f21686e6d726e736f6c7954550a6d20",
        INIT_38 => X"776e2072206d20454a0d6899613f748068454e0d65647420767420610d6f6920",
        INIT_39 => X"22652020206774687920e2206f2e616f20550a654a6e696c20226c6965646566",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000006979",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
         CLK     => clock,
         ADDR    => address,
         EN      => '1',
         WE      => we1,
         DI      => d_in_mem1,
         DIP     => "0",
         DO      => data_out(15 downto 8),
         SSR     => '0'
         );

   ----------------------------------------------------------------------------------
   -- bytes 7 a 0
   ----------------------------------------------------------------------------------
    block_0: RAMB16_S9
         generic map (
        INIT_00 => X"70207420747365574d5620490a737068206f6d6e6e650d206331410d6c646f52",
        INIT_01 => X"726e6961696c206e2067684149534f0a3f6374207265726e2066203f6161746f",
        INIT_02 => X"75650d6d2c6f746a7469614e4e45530a2e68756174207465777920206e736e6f",
        INIT_03 => X"72612074726f686565652074616e65686d2069206520686f0d61656f6f2c6f63",
        INIT_04 => X"6f656361666b202020475254460d612c2020475244540d7020206820656e6573",
        INIT_05 => X"732021626c682e20686e72656f6320475244540d626365656e72746f6e6f650a",
        INIT_06 => X"656565647375686c64656868616c43740a2e696520546c650a76726f686e6577",
        INIT_07 => X"20676e732068767420642e6565656c0d550a22654d680d20206c656f63206d6f",
        INIT_08 => X"650d6e206161653f6174656f6c0d2020687765726d200a6f6820626b20777268",
        INIT_09 => X"6c202069207761205461686565206e6c676d653f0a79656d4920726820656ce2",
        INIT_0A => X"656c65750d6f69e26e73806520992e656477205372737920666e6c6765680a65",
        INIT_0B => X"2c69720d6c202066416f65206120610a6564686e7920752e7073636d6d2e6565",
        INIT_0C => X"6520706f656c732072200a746f6e67207274726568756e2c73616872642c6175",
        INIT_0D => X"6f7365736e80696f6f2e6469646f61722020200a656169636f742c2073612065",
        INIT_0E => X"69e2636f6f69e261740a4c430d6179687920e220555354500d6b206965496165",
        INIT_0F => X"686e73796e2020666f2c7720796973737420436f65206c70656573540a636f6f",
        INIT_10 => X"656f6c54500d7968697348722c6c6973487273806520990d555354500d646177",
        INIT_11 => X"666420207268206861737920576e6e6520204f0a677220207774736e730d686d",
        INIT_12 => X"20756e6573730a68627574687474616820200d4f0a697477204149530d67206e",
        INIT_13 => X"65206e206853722020616f6572682020610d7273707461206563610a67666520",
        INIT_14 => X"676320416e20657068746ce2652073200a77206c20208079206e737363696e6f",
        INIT_15 => X"6773207475207473996e720d672c7273206e69767468200a6e65206473206d72",
        INIT_16 => X"686f657374722c572e7867206265722068462e614d656c736320202c544c540d",
        INIT_17 => X"65696b730a696d206f6e6320202c0a746520206e7361656f65206e6169656f65",
        INIT_18 => X"65722c614d73692c6e54590a73796f656557616977772c0a4c430d7374746c49",
        INIT_19 => X"73804c540d206f52750d550a2e6969796d736f206354742065207473616e6c41",
        INIT_1A => X"61746e2c65656c7065202065486561684c6f6c6765746e0d550a2e6f6969612c",
        INIT_1B => X"7969656e207461206165727464770d7564652d77616f69206f6d666720722c72",
        INIT_1C => X"72206f0d6572686969652c7720742e206520652065702066682e6d7269696475",
        INIT_1D => X"0d6561206c20636e20660a410a2e65202061656e652d200d77206866756e6365",
        INIT_1E => X"3f2065207365490a742061656120626d67610d72652068484c430d6875202080",
        INIT_1F => X"6f702d63746c200a7467206d6e6d652080596c206420686f6d656e6f6c750d20",
        INIT_20 => X"690d652074202e206120200a74202054500d6573738065756854590a61686299",
        INIT_21 => X"69616159746820616c0d6520992c6165726e74200a617720756563746e202072",
        INIT_22 => X"63740d420d73656d6c68742069756520800d61722169722c69722e2c75426f78",
        INIT_23 => X"6e75696875776820770d69726e6620686962746579650a696d6c206c20777265",
        INIT_24 => X"752077617066206199654a69224d0d2e78482e6765e262207620656765770d61",
        INIT_25 => X"6f6720746f200d74642069696e756f2c6c0a6973696c67746e736f690d686572",
        INIT_26 => X"73467320737369656c6e6857682020686f6e20752c672047454a0d6965746820",
        INIT_27 => X"642c6c6e202048450a2e6be26d20682070207041687420618069696173686174",
        INIT_28 => X"6e7420732020697220680a4d0d72726975756574206c69697954550a6f72616c",
        INIT_29 => X"520d6180657066616868652020736154550a6965747574206c6f746761790a64",
        INIT_2A => X"490a2e7273696d6e202c6c206668226873200a6b496520e261796c20206d684f",
        INIT_2B => X"20616e796d6921726c7773654f70796f6e0d4f0a6f6520746869687079766e0a",
        INIT_2C => X"2077736d6922756820777372656d6f6d4d530a2e62e279737554550a72736948",
        INIT_2D => X"642c6c6f200a732020792020726f652c65627220550a656d682057450a226820",
        INIT_2E => X"6868766c53656f6f61616165756c202e7464616f617267202072497374202077",
        INIT_2F => X"6f20774f560a2e648066206520216f20640d6c43657322734f520d7765207573",
        INIT_30 => X"65206f6f72726e6c676154500d746e6d206d546149200a4d0d74202073722020",
        INIT_31 => X"6f2e656573686f6e202e2020682068686f6565200d646f6561736f6e69616157",
        INIT_32 => X"756c0d656d20800d6165202c2079686968206220e220686f6f652063204d2e69",
        INIT_33 => X"2020722020200a520d6e6c676f6968656e65686f54550a74206e627265647475",
        INIT_34 => X"6854550a6972206f626e207420720d550a6f66756e2077742073740a490a2e65",
        INIT_35 => X"726568206f73202061697347454a0d6e6e20550a6320206f612c686f66686880",
        INIT_36 => X"676f6f736e682c614d642c6f69616920697420550a656e656d20652065670aa8",
        INIT_37 => X"2068626f640a746f6e6b61776e6579655465206f206675206c6e4d454a0d6574",
        INIT_38 => X"6f656461497941490a3f7480687320e257530a2e6ea861616f73496865742065",
        INIT_39 => X"0a6e656c736e73546173742c436e206e454e0d692069776c650a617763206e4f",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000227865",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
         CLK     => clock,
         ADDR    => address,
         EN      => '1',
         WE      => we0,
         DI      => d_in_mem0,
         DIP     => "0",
         DO      => data_out(7 downto 0),
         SSR     => '0'
         );

end data_mem_mod1;
